module alu_decoder(ALUOp, func3, op_5, func7_5, ALUControl);

    input[1:0] ALUOp;
    input[2:0] func3;
    input op_5,func7_5;
    wire[1:0] cont;
    output[2:0] ALUControl;

    assign cont = {op_5 , func7_5};

    assign ALUControl = (ALUOp == 2'b00) ? 3'b000 :
                        (ALUOp == 2'b01) ? 3'b001 :
                        ((ALUOp == 2'b10) & (func3 == 3'b000) & (cont == 2'b11))? 3'b001 :
                        ((ALUOp == 2'b10) & (func3 == 3'b000) & (cont != 2'b11))? 3'b000 :
                        ((ALUOp == 2'b10) & (func3 == 3'b010)) ? 3'b101 :
                        ((ALUOp == 2'b10) & (func3 == 3'b110)) ? 3'b011 :
                        ((ALUOp == 2'b10) & (func3 == 3'b111)) ? 3'b010 : 3'b000;

endmodule